`timescale 1ns / 1ps

module testbench();
    reg clk, rst;
    reg ready;
    reg[31:0] op1, op2;
    wire[31:0] res;
    wire done;
    parameter PERIOD = 12;
    parameter NUM_TEST = 20;
    reg [31:0] mem [0:NUM_TEST*3-1]; 
    integer i;


double_multiplier dut(
    .clk (clk),
    .rst (rst),
    .ready (ready),
    .op1 (op1),
    .op2 (op2),
    .res (res),
    .done (done)
);


initial begin   
    // Test 1
    mem[0] = 32'b00000000000000000000000000000000; //0.0
    mem[1] = 32'b11111111100000000000000000000000; //-inf
    mem[2] = 32'b11111111110000000000000000000000; //nan quiet
    
    // Test 2
    mem[3] = 32'b01111111100000000000000000000000; //+inf
    mem[4] = 32'b00000000000000000000000000000000; //0.0
    mem[5] = 32'b11111111110000000000000000000000; //nan quiet
    
    // Test 3
    mem[6] = 32'b01111111100000000000000000000110; //nan signal
    mem[7] = 32'b00111111101000000000000000000000; //1.25
    mem[8] = 32'b01111111100000000000000000000110; //nan signal
    
    // Test 4
    mem[9] = 32'b00111111101000000000000000000000; //1.25
    mem[10] = 32'b11111111100000000000010000000110; //nan signal
    mem[11] = 32'b11111111100000000000010000000110; //nan signal
    
    // Test 5
    mem[12] = 32'b00111111101000000000000000000000; //1.25
    mem[13] = 32'b00000000000000000000000000000000; //0.0
    mem[14] = 32'b00000000000000000000000000000000; //0.0
    
    // Test 6
    mem[15] = 32'b10000000000000000000000000000000; //-0.0
    mem[16] = 32'b00111111101000000000000000000000; //1.25
    mem[17] = 32'b10000000000000000000000000000000; //-0.0
    
    // Test 7
    mem[18] = 32'b11111111100000000000000000000000; //-inf
    mem[19] = 32'b01000000000000000000000000000000; //2.0
    mem[20] = 32'b11111111100000000000000000000000; //-inf
    
    // Test 8
    mem[21] = 32'b01000000000000000000000000000000; //2.0
    mem[22] = 32'b01111111100000000000000000000000; //inf
    mem[23] = 32'b01111111100000000000000000000000; //inf
    
    // Test 9
    mem[24] = 32'b00000000010000000000000000000000; //5.87747175411e-39 (DENOM)
    mem[25] = 32'b00000000010000000000000000000000; //5.87747175411e-39 (DENOM)
    mem[26] = 32'b00000000000000000000000000000000; //0.0
    
    // Test 10
    mem[27] = 32'b00111111110000000000000000000000; //1.5
    mem[28] = 32'b00000000010000000000000000000000; //5.87747175411e-39 (DENOM)
    mem[29] = 32'b00000000011000000000000000000000; //8.81620763117e-39 (DENOM)
    
    // Test 11
    mem[30] = 32'b00000000010000000000000000000000; //5.87747175411e-39 (DENOM)
    mem[31] = 32'b00111110110000000000000000000000; //0.375
    mem[32] = 32'b00000000000110000000000000000000; //2.20405190779e-39 (DENOM)
    
    // Test 12
    mem[33] = 32'b01100000000000000000000000000000; //36893488147419103232
    mem[34] = 32'b01100000000000000000000000000000; //36893488147419103232
    mem[35] = 32'b01111111100000000000000000000000; //+inf
    
    // Test 13
    mem[36] = 32'b01000010111101110111100011110010; //123.7362213134765625
    mem[37] = 32'b00111010101000010011011111110100; //0.0012300000526010990142822265625
    mem[38] = 32'b00111110000110111101100100100111; //0.15219555795192718505859375
    
    // Test 14
    mem[39] = 32'b01000010100100011100110011001101; //72.90000152587890625
    mem[40] = 32'b01000001000100000000000000000000; //9.0
    mem[41] = 32'b01000100001001000000011001100111; //656.10003662109375
    
    // Test 15
    mem[42] = 32'b01000000011111111111111111111110; //3.999999523162841796875
    mem[43] = 32'b01000000000000000000000000000001; //2.0000002384185791015625
    mem[44] = 32'b01000001000000000000000000000000; //8.0
    
    // Test 16
    mem[45] = 32'b01000001000000000000000000000000; //8.0
    mem[46] = 32'b00000000000000000000000000000001; //1.40129846432e-45 (DENOM)
    mem[47] = 32'b00000000000000000000000000001000; //1.12103877146e-44 (DENOM)
    
    // Test 17
    mem[48] = 32'b01000001100000000000000000000000; //16.0
    mem[49] = 32'b00000000010000000000000000000000; //5.87747175411e-39 (DENOM)
    mem[50] = 32'b00000010000000000000000000000000; //9.40395480658e-38
         
    // Test 18
    mem[51] = 32'b00111100000000000000000000000000; //0.0078125
    mem[52] = 32'b00000011100000000000000000000000; //7.52316384526e-37
    mem[53] = 32'b00000000010000000000000000000000; //5.87747175411e-39 (DENORM) 
    
    // Test 19
    mem[54] = 32'b01000001010110000000000000000000; //13.5
    mem[55] = 32'b00111111100000000000000000000000; //1.0
    mem[56] = 32'b01000001010110000000000000000000; //13.5
         
    // Test 20
    mem[57] = 32'b01000000000000000000000000000000; //2.0
    mem[58] = 32'b01000000001000000000000000000000; //2.5
    mem[59] = 32'b01000000101000000000000000000000; //5.0 
end


always #(PERIOD/2) clk  <= !clk; // Set clock

initial 
begin    
    // Init
    clk <= 1'b1;
    ready <= 1'b0;
    rst <= 1'b0;
    
    // Wait for startup FPGA
    #(PERIOD*20);
    
    // Reset
    #PERIOD;
    rst <= 1'b1;
    #PERIOD;
    rst <= 1'b0;    
    
    // Test: Verilog vs VHDL
    $display("###############");
    $display("VERILOG vs VHDL");
    i = 0;
    while (i < NUM_TEST * 3) begin  
        #(PERIOD/2);      
        #PERIOD;
        ready <= 1'b1;
        #PERIOD;
        ready <= 1'b0;
        op1 <= mem[i];
        op2 <= mem[i+1];
        #PERIOD;
        #PERIOD;
        @(posedge done) #(PERIOD/2);
        if (res == mem[i+2])
            $display("TEST VERILOG %d OK", 1+i/3);
        else
            $display("TEST VERILOG %d FAILED -> res= %b -> correct= %b", 1+i/3, res, mem[i+2]);
        #PERIOD;
        if (res == mem[i+2])
            $display("TEST VHDL    %d OK", 1+i/3);
        else
            $display("TEST VHDL    %d FAILED -> res= %b -> correct= %b", 1+i/3, res, mem[i+2]);    
        #(PERIOD/2);    
        i = i + 3;
    end    
    
    // Test: Verilog and VHDL
    $display("###############");
    $display("VERILOG and VHDL");
    i = 0;
    while (i < NUM_TEST * 3) begin 
        #(PERIOD/2);       
        #PERIOD;
        ready <= 1'b1;
        #PERIOD;
        ready <= 1'b0;
        op1 <= mem[i];
        op2 <= mem[i+1];
        #PERIOD;
        op1 <= mem[i+3];
        op2 <= mem[i+4];
        #PERIOD;
        @(posedge done) #(PERIOD/2);
        if (res == mem[i+2])
            $display("TEST VERILOG %d OK", 1+i/3);
        else
            $display("TEST VERILOG %d FAILED -> res= %b", 1+i/3, res);
        #PERIOD;
        if (res == mem[i+5])
            $display("TEST VHDL    %d OK", 2+i/3);
        else
            $display("TEST VHDL    %d FAILED -> res= %b", 2+i/3, res);  
        #(PERIOD/2);      
        i = i + 6;
    end
end


endmodule
