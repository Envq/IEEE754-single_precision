`timescale 1ns / 1ps

module testbench();
    reg clk, rst;
    reg ready;
    reg[31:0] op1, op2;
    wire[31:0] res;
    wire done;
    parameter PERIOD = 10;//7.598;
    parameter SIZE_TEST = 10;
    reg [31:0] mem [0:SIZE_TEST*3-1]; 
    integer i;


double_multipler top_level(
    .clk (clk),
    .rst (rst),
    .ready (ready),
    .op1 (op1),
    .op2 (op2),
    .res (res),
    .done (done)
);


initial begin
    //Test1
    mem[0] = 32'b11111111100000000000000000000000; //-inf
    mem[1] = 32'b01000000000000000000000000000000; //2.0
    mem[2] = 32'b11111111100000000000000000000000; //-inf
    
    //Test2
    mem[3] = 32'b00111111101000000000000000000000; //1.25
    mem[4] = 32'b00000000000000000000000000000000; //0.0
    mem[5] = 32'b00000000000000000000000000000000; //0.0
    
    //Test3
    mem[6] = 32'b11111111100000000000000000000000; //-inf
    mem[7] = 32'b00000000000000000000000000000000; //0.0
    mem[8] = 32'b11111111111111111111111111111111; //-nan
    
    //Test4
    mem[9] = 32'b01111111100000000000000000000000; //+inf
    mem[10] = 32'b00000000000000000000000000000000; //0.0
    mem[11] = 32'b01111111111111111111111111111111; //+nan
    
    //Test5
    mem[12] = 32'b01000001100000100000000000000000; //16.25
    mem[13] = 32'b01000001000100000000000000000000; //9.0
    mem[14] = 32'b01000011000100100100000000000000; //146.25
    
    //Test6
    mem[15] = 32'b01000001101100000000000000000000; //22.0
    mem[16] = 32'b11000000101000000000000000000000; //-5.0
    mem[17] = 32'b11000010110111000000000000000000; //-110.0
    
    //Test7 //1|011 even
    mem[18] = 32'b01000000010110011001100110011010; //3.400000095367431640625
    mem[19] = 32'b01000000010110011001100110011010; //3.400000095367431640625
    mem[20] = 32'b01000001001110001111010111000011; //11.56000041961669921875
    
    //Test8 //1|111 even+inf
    mem[21] = 32'b01000010101001111010100011110110; //83.8300018310546875
    mem[22] = 32'b00111110000011110101110000101001; //0.14000000059604644775390625
    mem[23] = 32'b01000001001110111100011101111010; //11.7362003326416015625
    
    //Test9 //100 even+inf
    mem[24] = 32'b01000010111101110111100011110010; //123.7362213134765625
    mem[25] = 32'b00111010101000010011011111110100; //0.0012300000526010990142822265625
    mem[26] = 32'b00111110000110111101100100100111; //0.15219555795192718505859375
    
    //Test10  //010 inf
    mem[27] = 32'b01000010100100011100110011001101; //72.90000152587890625
    mem[28] = 32'b01000001000100000000000000000000; //9.0
    mem[29] = 32'b01000100001001000000011001100111; //656.10003662109375
    
    //Test10 //110 even+inf
    //mem[27] = 32'b01001001011101000010010000000000; //1000000.0
    //mem[28] = 32'b01001001010110010000001110001110; //888888.875
    //mem[29] = 32'b01010011010011101111010111101000; //888888885248
    
    //Test12 VHDL
    //mem[33] = 32'b01000010100100011100110011001101; //72.9
    //mem[34] = 32'b01000001000100000000000000000000; //9.0
    //mem[35] = 32'b01000100001001000000011001100110; //656.1
end

       

always #(PERIOD/2) clk  <= !clk; // Set clock
initial 
begin
    //Init
    clk <= 1'b1;
    ready <= 1'b0;
    rst <= 1'b0;
    i <= 0;
    
    // Reset
    #PERIOD;
    rst <= 1'b1;
    #PERIOD;
    rst <= 1'b0;
    
    
        // Test
    while (i < SIZE_TEST * 3) begin        
        #PERIOD;
        ready <= 1'b1;
        op1 <= mem[i];
        op2 <= mem[i+1];
        #PERIOD;
        op1 <= mem[i+3];
        op2 <= mem[i+4];
        #PERIOD;
        ready <= 1'b0;
        @(posedge done) #PERIOD;
        if (res == mem[i+2])
            $display("TEST VERILOG %d OK", 1+i/3);
        else
            $display("TEST VERILOG %d FAILED -> res= %b", 1+i/3, res);
        #PERIOD;
        if (res == mem[i+5])
            $display("TEST VHDL    %d OK", 2+i/3);
        else
            $display("TEST VHDL    %d FAILED -> res= %b", 2+i/3, res);        
        i = i + 6;
    end

end



endmodule
